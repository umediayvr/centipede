<?xml version="1.0" encoding="UTF-8"?>
<ColorDecisionList xmlns="urn:ASC:CDL:v1.01">
	<ColorDecision>
		<ColorCorrection id="034_SCR_030_cdl">
			<Error>saturation missing or malformed - using identity</Error>
			<SOPNode>
				<Slope>1.1 1.2 1.3</Slope>
				<Offset>0.1 0.2 0.3</Offset>
				<Power>1.4 1.5 1.6</Power>
			</SOPNode>
			<SatNode>
				<Saturation>1</Saturation>
			</SatNode>
		</ColorCorrection>
	</ColorDecision>
</ColorDecisionList>
